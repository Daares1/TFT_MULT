--------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.Std_Logic_1164.all;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
ENTITY Configurable_U2 IS
  PORT(
      O0 : OUT std_logic;
      O1 : OUT std_logic;
      O2 : OUT std_logic;
      O3 : OUT std_logic;
      O4 : OUT std_logic;
      I : IN std_logic_vector(4 downto 0)
  );
END Configurable_U2;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
ARCHITECTURE structure OF Configurable_U2 IS
BEGIN
    O0 <= I(0);
    O1 <= I(1);
    O2 <= I(2);
    O3 <= I(3);
    O4 <= I(4);
END structure;
--------------------------------------------------------------------------------
