--------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.Std_Logic_1164.all;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
ENTITY Configurable_U3 IS
  PORT(
      I0 : IN std_logic;
      I1 : IN std_logic;
      I2 : IN std_logic;
      I3 : IN std_logic;
      I4 : IN std_logic;
      I5 : IN std_logic;
      I6 : IN std_logic;
      I7 : IN std_logic;
      O : OUT std_logic_vector(7 downto 0)
  );
END Configurable_U3;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
ARCHITECTURE structure OF Configurable_U3 IS
BEGIN
    O(0) <= I0;
    O(1) <= I1;
    O(2) <= I2;
    O(3) <= I3;
    O(4) <= I4;
    O(5) <= I5;
    O(6) <= I6;
    O(7) <= I7;
END structure;
--------------------------------------------------------------------------------
